module regs (
    input logic[4:0] read_reg_1,
    input logic[4:0] read_reg_2,
    input logic[4:0] write_reg,
    input logic[31:0] write_data,
    output logic[31:0] read_data_1,
    output logic[31:0] read_data_2
);
    
endmodule