module alu (
    input logic[31:0] data_1,
    input logic[31:0] data_2,
    input logic[5:0] fn,
    output logic[31:0] r,
    output logic zero
);
    
endmodule